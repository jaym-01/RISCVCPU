module top(
    input logic clk,
    input logic rst,
    output logic [31:0] a0;
);



endmodule
