module top #(
    parameter A_WIDTH = 20,
    parameter D_WIDTH = 32
) (
    input logic clk, 
);
    
endmodule